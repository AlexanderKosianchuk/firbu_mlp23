library verilog;
use verilog.vl_types.all;
entity sdInitTest is
end sdInitTest;
