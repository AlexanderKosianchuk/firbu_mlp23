library verilog;
use verilog.vl_types.all;
entity PeriphUSBTest is
end PeriphUSBTest;
