library verilog;
use verilog.vl_types.all;
entity sdTest is
end sdTest;
