library verilog;
use verilog.vl_types.all;
entity movingAverageTest is
end movingAverageTest;
