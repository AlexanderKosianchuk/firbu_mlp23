library verilog;
use verilog.vl_types.all;
entity FATupdeterTest is
end FATupdeterTest;
